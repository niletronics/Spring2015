module fsm(ten,twenty,ready,dispense,returnten,bill);

input ten,twenty;
output ready,dispense,returnten,bill;



