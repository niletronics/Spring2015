module leadadder_tb();
parameter width = 4;
reg [width-1:0] InA, InB;
reg InC;
